----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
----------------------------------------------------------------------------------
ENTITY RP_top IS
  PORT(
    BTN             : IN  STD_LOGIC_VECTOR (3 DOWNTO 0);
    SW              : IN  STD_LOGIC_VECTOR (3 DOWNTO 0);
    LED             : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
  );
END RP_top;
----------------------------------------------------------------------------------
ARCHITECTURE Structural OF RP_top IS
----------------------------------------------------------------------------------



----------------------------------------------------------------------------------
BEGIN
----------------------------------------------------------------------------------


----------------------------------------------------------------------------------
END Structural;
----------------------------------------------------------------------------------
